library verilog;
use verilog.vl_types.all;
entity risc_cpu_tb is
end risc_cpu_tb;
