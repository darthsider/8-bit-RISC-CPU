library verilog;
use verilog.vl_types.all;
entity program_counter is
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        \in\            : in     vl_logic_vector(7 downto 0);
        load            : in     vl_logic;
        inc             : in     vl_logic;
        \out\           : out    vl_logic_vector(7 downto 0)
    );
end program_counter;
