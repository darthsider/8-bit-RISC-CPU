library verilog;
use verilog.vl_types.all;
entity tb_proRISC is
end tb_proRISC;
